 //------------------------------------------------------------------------------
 // Project      : ALU 
 // File Name    : alu_sequencer.sv
 // Developers   : T5
 // Created Date : 2024
 // Version      : V1.0
 //------------------------------------------------------------------------------
 // Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
 //------------------------------------------------------------------------------
 
class alu_sequencer extends uvm_component;
    `uvm_uvm_component_utils(alu_sequencer)

    function new(string name = "alu_sequencer");
        super.new(name);
    endfunction

    // Additional implementation details for uvm_component go here

endclass
