 //------------------------------------------------------------------------------
 // Project      : ALU 
 // File Name    : alu_sequence_item.sv
 // Developers   : T5
 // Created Date : 2024
 // Version      : V1.0
 //------------------------------------------------------------------------------
 // Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
 //------------------------------------------------------------------------------
 
class alu_sequence_item extends uvm_object;
    `uvm_uvm_object_utils(alu_sequence_item)

    function new(string name = "alu_sequence_item");
        super.new(name);
    endfunction

    // Additional implementation details for uvm_object go here

endclass
