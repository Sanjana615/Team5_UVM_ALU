 //------------------------------------------------------------------------------
 // Project      : ALU 
 // File Name    : alu_test.sv
 // Developers   : T5
 // Created Date : 2024
 // Version      : V1.0
 //------------------------------------------------------------------------------
 // Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
 //------------------------------------------------------------------------------
 
class alu_test extends uvm_component;
    `uvm_uvm_component_utils(alu_test)

    function new(string name = "alu_test");
        super.new(name);
    endfunction

    // Additional implementation details for uvm_component go here

endclass
